module rjsc5(
  input clk,
  input reset
);

endmodule